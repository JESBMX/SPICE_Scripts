A3_E2_BJT_Curves_Tracer
* -------------------------------------------
*      A3_E2 - BJT Curves Tracer

* BJT Under Test
* Q1	c	b	0	Q2N2222
* Q1	c	b	0	Q2N2222A
Q1	c	b	0	Q2N3904

* Sources definition
Vce	c	0	DC	1V
Ib	0	bx	DC	1uA
Vb	b	bx	DC	0V

* Models
.MODEL Q2N2222 NPN
	+ (IS=3.108E-15 XTI=3 EG=1.11 VAF=131.5 BF=217.5
	+ NE=1.541 ISE=190.7E-15 IKF=1.296 XTB=1.5 BR=6.18
	+ NC=2 ISC=0 IKR=0 RC=1 CJC=14.57E-12 VJC=.75
	+ MJC=.3333 FC=.5 CJE=26.08E-12 VJE=.75 MJE=.3333
	+ TR=51.35E-9 TF=451E-12 ITF=.1 VTF=10 XTF=2)

.MODEL Q2N2222A NPN
	+ IS=3.88184e-14 BF=929.846 NF=1.10496 VAF=16.5003
	+ IKF=0.019539 ISE=1.0168e-11 NE=1.94752 BR=48.4545
	+ NR=1.07004 VAR=40.538 IKR=0.19539 ISC=1.0168e-11
	+ NC=4 RB=0.1 IRB=0.1 RBM=0.1
	+ RE=0.0001 RC=0.426673 XTB=0.1 XTI=1
	+ EG=1.05 CJE=2.23677e-11 VJE=0.582701 MJE=0.63466
	+ TF=4.06711e-10 XTF=3.92912 VTF=17712.6 ITF=0.4334
	+ CJC=2.23943e-11 VJC=0.576146 MJC=0.632796 XCJC=1
	+ FC=0.170253 CJS=0 VJS=0.75 MJS=0.5
	+ TR=1e-07 PTF=0 KF=0 AF=1

.MODEL Q2N3904 NPN
	+ IS=1.26532e-10 BF=206.302 NF=1.5 VAF=1000
	+ IKF=0.0272221 ISE=2.30771e-09 NE=3.31052 BR=20.6302
	+ NR=2.89609 VAR=9.39809 IKR=0.272221 ISC=2.30771e-09
	+ NC=1.9876 RB=5.8376 IRB=50.3624 RBM=0.634251
	+ RE=0.0001 RC=2.65711 XTB=0.1 XTI=1
	+ EG=1.05 CJE=4.64214e-12 VJE=0.4 MJE=0.256227
	+ TF=4.19578e-10 XTF=0.906167 VTF=8.75418 ITF=0.0105823
	+ CJC=3.76961e-12 VJC=0.4 MJC=0.238109 XCJC=0.8
	+ FC=0.512134 CJS=0 VJS=0.75 MJS=0.5
	+ TR=6.82023e-08 PTF=0 KF=0 AF=1

* Analysis definition
.control
destroy all

* DC Vce 0V 30V 0.1V Ib 0.5uA 300uA 50uA
* Ic = -i(Vce)
* PLOT Ic xlabel Vce ylabel Ic

DC Ib 0.5uA 300uA 5uA Vce 1V 28V 9V
beta = i(Vce)/i(Vb)
PLOT beta xunits A yunits b xlabel Ib ylabel Beta
.endc

.end