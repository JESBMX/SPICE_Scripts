Series_Clipper
* -----------------------------------------------------
*                    Series Clipper

Vs   in  0     DC 0V   AC 1V   SIN(0V 4V 1KHz)
Rs   in  in2   1
*D1   in2 out   D1N4004
D1   in2 out   ideal_diode
VR   out out2  DC  2V
RL   out2 0    100

* 1N4004 - 1A 400V General Purpose Rectifier
* Fairchild (now National Semiconductors)
.MODEL  D1N4004  D (IS=3.699E-09 RS=1.756E-02 N=1.774
+       XTI=3.0 EG=1.110 CJO=1.732E-11 M=0.3353
+       VJ=0.3905 FC=0.5 BV=400 IBV=1.0E-03)

* Quasi Ideal Diode
.model ideal_diode D (Is=1pA n=0.01)

*.TRAN 10E-6 4E-3
*.plot tran v(in) v(out)
*.end

.control
TRAN 10E-6 4E-3
PLOT v(in) v(out)
.endc

.end